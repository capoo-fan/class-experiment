module top (
    input wire clk,        // 100MHz ʱ��
    input wire S1,          // �첽��λ
    input wire S3,          // ���Ͱ���
    input wire uart_rx,    // UART ����
    input wire SW0,        // ���� SW0,string_match �ͷ���ѧ�ŵ��л��ź�
    output wire uart_tx,   // UART ����
    output wire [7:0] led_en,  // �����λѡ
    output wire [7:0] led_cx   // ����ܶ�ѡ
  );

  wire rst = S1;

  // S3
  wire s3_debounced;
  wire s3_posedge;

  // UART ����
  wire recv_valid;
  wire [7:0] recv_data;

  // �������ʾ
  wire [39:0] display_data; // ���ӵ� led_ctrl_unit ������


  wire s3_mode_tx;      //send mode
  wire match_mode_tx; //string match mode

  assign uart_tx = (SW0 == 1'b0) ? s3_mode_tx : match_mode_tx;

  // ���� S3 ����
  debounce #(
             .cnt_max(2_000_000)
           ) u_debounce_s3 (
             .clk(clk),
             .rst(rst),
             .button_in(S3),
             .button_out(s3_debounced)
           );

  // S3 �����ؼ��
  edge_detect u_edge_detect_s3 (
                .clk(clk),
                .rst(rst),
                .signal(s3_debounced),
                .pos_edge(s3_posedge)
              );

  // UART ����
  uart_recv u_uart_recv (
              .clk(clk),
              .rst(rst),
              .din(uart_rx),
              .valid(recv_valid),
              .data(recv_data)
            );

  // UART ����������ʾ�߼�
  // ��������յ������ݲ�����39λ��ʾ����
  display_logic u_display_logic (
                  .clk(clk),
                  .rst(rst),
                  .valid(recv_valid),
                  .recv_data(recv_data),
                  .display_data(display_data) // ����� led_ctrl
                );

  // 8 λ���������
  led_ctrl_unit #(
                  .time_max(100_000 - 1) // 1ms ˢ����
                ) u_led_ctrl (
                  .rst(rst),
                  .clk(clk),
                  .display(display_data), // ���ӵ� display_logic �����
                  .led_en(led_en),
                  .led_cx(led_cx)
                );

  send_ctrl u_send_ctrl (
              .clk(clk),
              .rst(rst),
              .s3(s3_posedge),
              .uart_tx(s3_mode_tx)
            );

  string_match u_string_match (
                 .clk(clk),
                 .rst(rst),
                  .valid(recv_valid),
                 .recv_data(recv_data),
                 .uart_tx(match_mode_tx)
               );

endmodule
