`timescale 1ns / 1ps
module tb_top;
  reg clk;
  reg S1;       // ��λ
  reg S2;       // ��ͣ
  reg S3;       // ����
  reg SW0;      // �ܿ���

  // ��Ӧ top ģ��� output
  wire [7:0] led_en;
  wire [7:0] led_cx;

  // �۲��������ʾ������
  wire [31:0] data_display;
  assign data_display = u_top.display;

  // ����
  top #(
        .clock_max(1000 - 1),  // 10us 30�μ���������
        .cnt_max(1000 ),   // 10us ����ʱ��
        .time_max(100-1)   // 1us ˢ��ʱ��
      )u_top (
        .clk(clk),
        .S1(S1),
        .S2(S2),
        .S3(S3),
        .SW0(SW0),
        .led_en(led_en),
        .led_cx(led_cx)
      );

  initial
    begin
      clk = 0;
    end
  always #5 clk = ~clk;

  initial
    begin
      S1 = 1;
      S2 = 0;
      S3 = 0;
      SW0 = 0; // ��ʼ״̬
      #10;

      S1=0;
      #10;
      // �ڲ����м�������ӦΪ 0

      SW0 = 1; // �����ܿ���

      // *** ��Ҫ��ʾ: ���·�˵�� (1) ***
      // 0.1s = 100,000,000 ns. ��������.
      // �ȴ� 3.5 �� 0.1s ����, �۲� DK1-DK0
      #(10000); // 10us ��, data_display[7:0] ӦΪ 8'h01
      #(10000); // 20us ��, data_display[7:0] ӦΪ 8'h02
      #(10000); // 30us ��, data_display[7:0] ӦΪ 8'h03

      // S2 ��ͣ
      S2 = 1;
      #(10000+1000);
      S2 = 0;

      // �ȴ� 2us, ����ֵ Ӧ�ñ����� 8'h03 ����
      #(20000);

      S2 = 1;
      #1000;
      S2 = 0; // �ٴΰ���, ģ��ë��

      #(10000); // 10us ��, ����ֵ���ɲ���


      // ���԰�����������
      S3 = 1;
      #10;
      S3 = 0; // ģ��ë��
      #10000;

      S3 = 1;
      #10;
      S3 = 0; // ģ��ë��
      #10000;

      S3 = 1;
      #10;
      S3 = 0; // ģ��ë��
      #10000;

      
      S3 = 1; // ��������
      #(10000+1000); // 10us ����ʱ��
      S3 = 0; // �ͷŰ���
      #(10000+1000);

      S3 = 1; 
      #(10000+1000); 
      S3 = 0; 
      #(10000+1000);

      // ��ʱ��������Ӧ��ֻ����������

      // (5) ���� SW0 �ر���ʾ
      SW0 = 0;
      #10000; // �ȴ� 10us����ʾȫ��
      $finish; 
    end

endmodule
